//develop control in parallel with datapath 
