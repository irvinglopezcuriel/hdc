//develop datapath in parallel with control 
