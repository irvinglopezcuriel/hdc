 // this is the encoding control file
